CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 570 30 120 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
244318226 0
0
6 Title:
5 Name:
0
0
0
63
13 Logic Switch~
5 138 706 0 1 11
0 3
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V15
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
45093.2 0
0
13 Logic Switch~
5 1485 443 0 1 11
0 10
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V14
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
45093.2 0
0
13 Logic Switch~
5 848 453 0 1 11
0 14
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V12
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3124 0 0
2
45093.2 0
0
13 Logic Switch~
5 852 364 0 1 11
0 16
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V11
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3421 0 0
2
45093.2 0
0
13 Logic Switch~
5 150 402 0 1 11
0 19
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8157 0 0
2
45093.2 1
0
13 Logic Switch~
5 1475 226 0 1 11
0 28
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5572 0 0
2
45093.2 0
0
13 Logic Switch~
5 1478 113 0 1 11
0 29
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8901 0 0
2
45093.2 0
0
13 Logic Switch~
5 699 113 0 1 11
0 33
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7361 0 0
2
45093.2 0
0
13 Logic Switch~
5 136 197 0 1 11
0 39
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4747 0 0
2
45093.2 0
0
13 Logic Switch~
5 143 84 0 1 11
0 40
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
972 0 0
2
45093.2 0
0
7 Ground~
168 468 776 0 1 3
0 2
0
0 0 53360 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3472 0 0
2
45093.2 0
0
12 Hex Display~
7 476 657 0 18 19
10 5 4 2 2 0 0 0 0 0
0 1 1 0 1 1 0 1 2
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP7
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
9998 0 0
2
45093.2 0
0
5 4027~
219 272 757 0 7 32
0 41 3 6 3 42 4 5
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U8B
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 8 0
1 U
3536 0 0
2
45093.2 4
0
7 Pulser~
4 195 744 0 10 12
0 43 44 6 45 0 0 10 10 3
8
0
0 0 4656 0
0
3 V16
-11 -28 10 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
4597 0 0
2
45093.2 3
0
14 Logic Display~
6 360 690 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L14
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3835 0 0
2
45093.2 2
0
14 Logic Display~
6 423 689 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L13
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3670 0 0
2
45093.2 1
0
7 Ground~
168 1814 513 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5616 0 0
2
45093.2 0
0
12 Hex Display~
7 1824 392 0 18 19
10 8 7 2 2 0 0 0 0 0
0 1 1 0 1 1 0 1 2
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP6
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
9323 0 0
2
45093.2 0
0
9 Inverter~
13 1487 516 0 2 22
0 10 9
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U2B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
317 0 0
2
45093.2 0
0
14 Logic Display~
6 1770 426 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L12
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3108 0 0
2
45093.2 0
0
14 Logic Display~
6 1707 427 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L11
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4299 0 0
2
45093.2 0
0
7 Pulser~
4 1542 481 0 10 12
0 46 47 11 48 0 0 10 10 3
8
0
0 0 4656 0
0
3 V13
-11 -28 10 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
9672 0 0
2
45093.2 0
0
5 4027~
219 1619 494 0 7 32
0 49 10 11 9 50 7 8
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U8A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 8 0
1 U
7876 0 0
2
45093.2 0
0
7 Ground~
168 1218 447 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
6369 0 0
2
45093.2 0
0
12 Hex Display~
7 1231 359 0 18 19
10 13 12 2 2 0 0 0 0 0
0 1 1 1 1 0 0 1 3
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP5
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
9172 0 0
2
45093.2 0
0
14 Logic Display~
6 1156 336 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L10
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7100 0 0
2
45093.2 0
0
14 Logic Display~
6 1083 340 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3820 0 0
2
45093.2 0
0
7 Pulser~
4 886 409 0 10 12
0 51 52 15 53 0 0 10 10 3
8
0
0 0 4656 0
0
2 V8
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
7678 0 0
2
45093.2 0
0
6 74112~
219 978 416 0 7 32
0 54 16 15 14 55 12 13
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U7A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 7 0
1 U
961 0 0
2
45093.2 0
0
5 7412~
219 275 403 0 4 22
0 18 19 22 21
0
0 0 624 0
4 7412
-7 -24 21 -16
3 U6A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 6 0
65 0 0 0 3 1 6 0
1 U
3178 0 0
2
45093.2 10
0
5 7412~
219 273 514 0 4 22
0 22 19 17 20
0
0 0 624 0
4 7412
-7 -24 21 -16
3 U4C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 6 0
65 0 0 0 3 3 4 0
1 U
3409 0 0
2
45093.2 9
0
10 2-In NAND~
219 387 410 0 3 22
0 21 17 18
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
3951 0 0
2
45093.2 8
0
10 2-In NAND~
219 387 506 0 3 22
0 18 20 17
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
8885 0 0
2
45093.2 7
0
14 Logic Display~
6 499 375 0 1 2
10 18
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3780 0 0
2
45093.2 6
0
14 Logic Display~
6 575 370 0 1 2
10 17
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9265 0 0
2
45093.2 5
0
7 Pulser~
4 136 448 0 10 12
0 56 57 22 58 0 0 10 10 3
8
0
0 0 4656 0
0
3 V10
-10 -28 11 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
9442 0 0
2
45093.2 4
0
12 Hex Display~
7 635 382 0 16 19
10 18 17 2 2 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP4
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
9424 0 0
2
45093.2 3
0
7 Ground~
168 625 485 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
9968 0 0
2
45093.2 2
0
7 Ground~
168 1953 196 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
9281 0 0
2
45093.2 0
0
12 Hex Display~
7 1963 93 0 16 19
10 26 25 2 2 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP3
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
8464 0 0
2
45093.2 0
0
7 Pulser~
4 1464 159 0 10 12
0 59 60 27 61 0 0 10 10 3
8
0
0 0 4656 0
0
2 V7
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
7168 0 0
2
45093.2 0
0
14 Logic Display~
6 1903 81 0 1 2
10 25
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3171 0 0
2
45093.2 0
0
14 Logic Display~
6 1827 86 0 1 2
10 26
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4139 0 0
2
45093.2 0
0
10 2-In NAND~
219 1715 217 0 3 22
0 26 23 25
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U3D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
6435 0 0
2
45093.2 0
0
10 2-In NAND~
219 1715 121 0 3 22
0 24 25 26
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
5283 0 0
2
45093.2 0
0
5 7412~
219 1601 225 0 4 22
0 27 28 26 23
0
0 0 624 0
4 7412
-7 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 6 0
65 0 0 0 3 2 4 0
1 U
6874 0 0
2
45093.2 0
0
5 7412~
219 1603 114 0 4 22
0 25 29 27 24
0
0 0 624 0
4 7412
-7 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 6 0
65 0 0 0 3 1 4 0
1 U
5305 0 0
2
45093.2 0
0
10 2-In NAND~
219 858 121 0 3 22
0 33 36 35
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
34 0 0
2
45093.2 10
0
10 2-In NAND~
219 857 230 0 3 22
0 36 32 34
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
969 0 0
2
45093.2 9
0
10 2-In NAND~
219 987 126 0 3 22
0 35 30 31
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U1D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
8402 0 0
2
45093.2 8
0
10 2-In NAND~
219 989 229 0 3 22
0 31 34 30
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
3751 0 0
2
45093.2 7
0
14 Logic Display~
6 1094 91 0 1 2
10 31
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4292 0 0
2
45093.2 6
0
14 Logic Display~
6 1166 87 0 1 2
10 30
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6118 0 0
2
45093.2 5
0
7 Pulser~
4 677 170 0 10 12
0 62 63 36 64 0 0 10 10 3
8
0
0 0 4656 0
0
2 V4
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
34 0 0
2
45093.2 4
0
9 Inverter~
13 743 241 0 2 22
0 33 32
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
6357 0 0
2
45093.2 3
0
12 Hex Display~
7 1227 101 0 18 19
10 31 30 2 2 0 0 0 0 0
0 1 1 0 1 1 0 1 2
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
319 0 0
2
45093.2 2
0
7 Ground~
168 1221 198 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3976 0 0
2
45093.2 1
0
7 Ground~
168 458 186 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7634 0 0
2
45093.2 0
0
12 Hex Display~
7 468 77 0 18 19
10 38 37 2 2 0 0 0 0 0
0 1 1 1 1 0 0 1 3
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
523 0 0
2
45093.2 0
0
14 Logic Display~
6 413 47 0 1 2
10 37
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6748 0 0
2
45093.2 0
0
14 Logic Display~
6 345 52 0 1 2
10 38
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6901 0 0
2
45093.2 0
0
10 2-In NAND~
219 241 202 0 3 22
0 38 39 37
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
842 0 0
2
45093.2 0
0
10 2-In NAND~
219 242 97 0 3 22
0 40 37 38
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3277 0 0
2
45093.2 0
0
85
0 1 2 0 0 4096 0 0 11 3 0 3
474 751
474 770
468 770
1 4 3 0 0 8320 0 1 13 0 0 4
150 706
150 776
248 776
248 739
3 4 2 0 0 8208 0 12 12 0 0 6
473 681
474 681
474 751
468 751
468 681
467 681
0 2 4 0 0 4112 0 0 12 6 0 4
422 739
480 739
480 681
479 681
0 1 5 0 0 4240 0 0 12 7 0 4
360 721
486 721
486 681
485 681
6 1 4 0 0 4240 0 13 16 0 0 3
302 739
423 739
423 707
7 1 5 0 0 16 0 13 15 0 0 3
296 721
360 721
360 708
3 3 6 0 0 4240 0 14 13 0 0 4
219 735
241 735
241 730
248 730
1 2 3 0 0 16 0 1 13 0 0 3
150 706
248 706
248 721
0 1 2 0 0 0 0 0 17 11 0 3
1817 488
1817 507
1814 507
3 4 2 0 0 4224 0 18 18 0 0 4
1821 416
1821 488
1815 488
1815 416
0 2 7 0 0 8192 0 0 18 14 0 3
1769 476
1827 476
1827 416
0 1 8 0 0 4224 0 0 18 15 0 3
1707 458
1833 458
1833 416
6 1 7 0 0 4224 0 23 20 0 0 3
1649 476
1770 476
1770 444
7 1 8 0 0 0 0 23 21 0 0 3
1643 458
1707 458
1707 445
2 4 9 0 0 8320 0 19 23 0 0 4
1490 534
1490 545
1595 545
1595 476
1 1 10 0 0 4096 0 2 19 0 0 4
1497 443
1497 483
1490 483
1490 498
3 3 11 0 0 4224 0 22 23 0 0 4
1566 472
1588 472
1588 467
1595 467
1 2 10 0 0 4224 0 2 23 0 0 3
1497 443
1595 443
1595 458
0 1 2 0 0 0 0 0 24 21 0 3
1224 428
1224 441
1218 441
3 4 2 0 0 0 0 25 25 0 0 4
1228 383
1228 428
1222 428
1222 383
0 2 12 0 0 8192 0 0 25 24 0 4
1155 398
1155 418
1234 418
1234 383
0 1 13 0 0 4224 0 0 25 25 0 5
1081 380
1170 380
1170 397
1240 397
1240 383
6 1 12 0 0 4224 0 29 26 0 0 3
1008 398
1156 398
1156 354
7 1 13 0 0 0 0 29 27 0 0 3
1002 380
1083 380
1083 358
1 4 14 0 0 4224 0 3 29 0 0 4
860 453
948 453
948 398
954 398
3 3 15 0 0 4224 0 28 29 0 0 4
910 400
933 400
933 389
948 389
1 2 16 0 0 4224 0 4 29 0 0 4
864 364
923 364
923 380
954 380
3 0 17 0 0 12416 0 31 0 0 40 5
249 523
228 523
228 538
483 538
483 506
1 0 18 0 0 12416 0 30 0 0 41 5
251 394
233 394
233 356
430 356
430 410
0 2 19 0 0 4224 0 0 31 44 0 3
194 402
194 514
249 514
4 2 20 0 0 8320 0 31 33 0 0 3
300 514
300 515
363 515
4 1 21 0 0 8320 0 30 32 0 0 3
302 403
302 401
363 401
0 1 2 0 0 0 0 0 38 35 0 3
627 457
625 457
625 479
3 4 2 0 0 0 0 37 37 0 0 4
632 406
632 457
626 457
626 406
0 2 17 0 0 0 0 0 37 40 0 3
575 450
638 450
638 406
0 1 18 0 0 0 0 0 37 41 0 4
495 410
495 427
644 427
644 406
1 0 18 0 0 0 0 33 0 0 41 5
363 497
347 497
347 471
458 471
458 410
2 0 17 0 0 0 0 32 0 0 40 5
363 419
335 419
335 458
443 458
443 506
3 1 17 0 0 0 0 33 35 0 0 3
414 506
575 506
575 388
3 1 18 0 0 0 0 32 34 0 0 3
414 410
499 410
499 393
3 0 22 0 0 4096 0 36 0 0 43 2
160 439
241 439
3 1 22 0 0 8320 0 30 31 0 0 4
251 412
241 412
241 505
249 505
1 2 19 0 0 0 0 5 30 0 0 4
162 402
243 402
243 403
251 403
4 2 23 0 0 8320 0 46 44 0 0 3
1628 225
1628 226
1691 226
4 1 24 0 0 8320 0 47 45 0 0 3
1630 114
1630 112
1691 112
0 1 2 0 0 0 0 0 39 48 0 3
1955 168
1953 168
1953 190
3 4 2 0 0 0 0 40 40 0 0 4
1960 117
1960 168
1954 168
1954 117
0 2 25 0 0 4096 0 0 40 55 0 3
1903 161
1966 161
1966 117
0 1 26 0 0 8192 0 0 40 56 0 4
1823 121
1823 138
1972 138
1972 117
3 0 26 0 0 12416 0 46 0 0 56 5
1577 234
1558 234
1558 257
1811 257
1811 121
1 0 25 0 0 12416 0 47 0 0 55 5
1579 105
1566 105
1566 52
1861 52
1861 217
1 0 26 0 0 0 0 44 0 0 56 5
1691 208
1675 208
1675 182
1786 182
1786 121
2 0 25 0 0 0 0 45 0 0 55 5
1691 130
1663 130
1663 169
1771 169
1771 217
3 1 25 0 0 0 0 44 42 0 0 3
1742 217
1903 217
1903 99
3 1 26 0 0 0 0 45 43 0 0 3
1742 121
1827 121
1827 104
3 0 27 0 0 4096 0 41 0 0 59 2
1488 150
1569 150
1 2 28 0 0 4224 0 6 46 0 0 4
1487 226
1569 226
1569 225
1577 225
3 1 27 0 0 8320 0 47 46 0 0 4
1579 123
1569 123
1569 216
1577 216
1 2 29 0 0 4224 0 7 47 0 0 4
1490 113
1571 113
1571 114
1579 114
0 1 2 0 0 0 0 0 57 62 0 3
1224 177
1224 192
1221 192
3 4 2 0 0 0 0 56 56 0 0 4
1224 125
1224 177
1218 177
1218 125
0 2 30 0 0 4096 0 0 56 70 0 3
1166 162
1230 162
1230 125
0 1 31 0 0 8320 0 0 56 71 0 4
1087 126
1087 146
1236 146
1236 125
2 2 32 0 0 4224 0 55 49 0 0 4
764 241
825 241
825 239
833 239
1 1 33 0 0 4224 0 8 55 0 0 3
711 113
711 241
728 241
1 1 33 0 0 0 0 8 48 0 0 3
711 113
711 112
834 112
1 0 31 0 0 0 0 51 0 0 71 5
965 220
951 220
951 192
1070 192
1070 126
2 0 30 0 0 12288 0 50 0 0 70 5
963 135
941 135
941 181
1051 181
1051 229
3 1 30 0 0 4224 0 51 53 0 0 3
1016 229
1166 229
1166 105
3 1 31 0 0 0 0 50 52 0 0 3
1014 126
1094 126
1094 109
3 2 34 0 0 4224 0 49 51 0 0 4
884 230
957 230
957 238
965 238
3 1 35 0 0 4224 0 48 50 0 0 4
885 121
955 121
955 117
963 117
3 0 36 0 0 4224 0 54 0 0 75 4
701 161
810 161
810 162
825 162
2 1 36 0 0 0 0 48 49 0 0 4
834 130
825 130
825 221
833 221
0 1 2 0 0 0 0 0 58 77 0 3
461 164
461 180
458 180
3 4 2 0 0 128 0 59 59 0 0 4
465 101
465 164
459 164
459 101
0 2 37 0 0 4096 0 0 59 84 0 3
413 143
471 143
471 101
0 1 38 0 0 8320 0 0 59 85 0 4
340 97
340 120
477 120
477 101
1 0 38 0 0 128 0 62 0 0 85 5
217 193
213 193
213 158
312 158
312 97
2 0 37 0 0 12288 0 63 0 0 84 5
218 106
204 106
204 150
298 150
298 202
1 2 39 0 0 4224 0 9 62 0 0 4
148 197
209 197
209 211
217 211
1 1 40 0 0 4224 0 10 63 0 0 4
155 84
210 84
210 88
218 88
3 1 37 0 0 4224 0 62 60 0 0 3
268 202
413 202
413 65
3 1 38 0 0 0 0 63 61 0 0 3
269 97
345 97
345 70
30
-19 0 0 0 400 0 0 0 0 0 0 0 23
12 Cooper Black
0 0 0 6
63 593 146 623
72 599 136 621
6 Task 7
-19 0 0 0 400 0 0 0 0 0 0 0 23
12 Cooper Black
0 0 0 1
81 659 109 689
88 666 101 688
1 T
-19 0 0 0 400 0 0 0 0 0 0 0 23
12 Cooper Black
0 0 0 6
1377 353 1462 383
1387 360 1451 382
6 Task 6
-19 0 0 0 400 0 0 0 0 0 0 0 23
12 Cooper Black
0 0 0 1
1435 411 1471 441
1445 418 1460 440
1 D
-19 0 0 0 400 0 0 0 0 0 0 0 23
12 Cooper Black
0 0 0 3
1532 504 1592 534
1541 511 1582 533
3 CLK
-19 0 0 0 400 0 0 0 0 0 0 0 23
12 Cooper Black
0 0 0 6
719 292 802 322
728 299 792 321
6 Task 5
-19 0 0 0 400 0 0 0 0 0 0 0 23
12 Cooper Black
0 0 0 1
804 435 835 465
813 442 825 464
1 J
-19 0 0 0 400 0 0 0 0 0 0 0 23
12 Cooper Black
0 0 0 3
801 380 861 410
810 387 851 409
3 CLK
-19 0 0 0 400 0 0 0 0 0 0 0 23
12 Cooper Black
0 0 0 1
808 341 840 371
817 348 830 370
1 S
-19 0 0 0 400 0 0 0 0 0 0 0 23
12 Cooper Black
0 0 0 1
91 369 119 399
98 376 111 398
1 T
-19 0 0 0 400 0 0 0 0 0 0 0 23
12 Cooper Black
0 0 0 6
40 317 123 347
49 323 113 345
6 Task 4
-19 0 0 0 400 0 0 0 0 0 0 0 23
12 Cooper Black
0 0 0 3
53 427 113 457
62 434 103 456
3 CLK
-19 0 0 0 400 0 0 0 0 0 0 0 23
12 Cooper Black
0 0 0 1
458 357 492 387
467 364 482 386
1 Q
-19 0 0 0 400 0 0 0 0 0 0 0 23
12 Cooper Black
0 0 0 2
533 357 571 387
542 363 561 385
2 Q'
-19 0 0 0 400 0 0 0 0 0 0 0 23
12 Cooper Black
0 0 0 6
1368 28 1453 58
1378 35 1442 57
6 Task 3
-19 0 0 0 400 0 0 0 0 0 0 0 23
12 Cooper Black
0 0 0 2
1861 68 1899 98
1870 74 1889 96
2 Q'
-19 0 0 0 400 0 0 0 0 0 0 0 23
12 Cooper Black
0 0 0 1
1786 68 1820 98
1795 75 1810 97
1 Q
-19 0 0 0 400 0 0 0 0 0 0 0 23
12 Cooper Black
0 0 0 1
1424 208 1459 238
1433 215 1449 237
1 K
-19 0 0 0 400 0 0 0 0 0 0 0 23
12 Cooper Black
0 0 0 3
1381 138 1441 168
1390 145 1431 167
3 CLK
-19 0 0 0 400 0 0 0 0 0 0 0 23
12 Cooper Black
0 0 0 1
1419 80 1452 110
1429 87 1441 109
1 J
-19 0 0 0 400 0 0 0 0 0 0 0 23
12 Cooper Black
0 0 0 6
641 31 724 61
650 38 714 60
6 Task 2
-19 0 0 0 400 0 0 0 0 0 0 0 23
12 Cooper Black
0 0 0 1
648 90 682 120
657 97 672 119
1 D
-19 0 0 0 400 0 0 0 0 0 0 0 23
12 Cooper Black
0 0 0 3
618 190 678 220
627 197 668 219
3 CLK
-19 0 0 0 400 0 0 0 0 0 0 0 23
12 Cooper Black
0 0 0 1
1050 63 1084 93
1059 70 1074 92
1 Q
-19 0 0 0 400 0 0 0 0 0 0 0 23
12 Cooper Black
0 0 0 2
1121 68 1161 98
1131 75 1150 97
2 Q'
-19 0 0 0 400 0 0 0 0 0 0 0 23
12 Cooper Black
0 0 0 6
29 15 112 45
38 22 102 44
6 Task 1
-19 0 0 0 400 0 0 0 0 0 0 0 23
12 Cooper Black
0 0 0 2
371 32 411 62
381 38 400 60
2 Q'
-19 0 0 0 400 0 0 0 0 0 0 0 23
12 Cooper Black
0 0 0 1
305 28 339 58
314 35 329 57
1 Q
-19 0 0 0 400 0 0 0 0 0 0 0 23
12 Cooper Black
0 0 0 1
89 172 123 202
98 179 113 201
1 R
-19 0 0 0 400 0 0 0 0 0 0 0 23
12 Cooper Black
0 0 0 1
93 58 125 88
102 65 115 87
1 S
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
